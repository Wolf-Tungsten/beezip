`define DEBUG_LOG

`ifdef DEBUG_LOG

// `define HASH_ENGINE_DEBUG_LOG

// `define MATCH_ENGINE_DEBUG_LOG

`ifdef MATCH_ENGINE_DEBUG_LOG

`define JOB_PE_DEBUG_LOG
`define MATCH_PE_DEBUG_LOG
`define SEQ_BUS_DEBUG_LOG
`define MESH_DEBUG_LOG

`endif // MATCH_ENGINE_DEBUG_LOG

`endif // DEBUG_LOG

`ifndef DATA_TYPES_V
`define DATA_TYPES_V

`include "parameters.v"

`endif DATA_TYPES_V
`ifndef UTIL_VH
`define UTIL_VH

`define TD #1

`endif